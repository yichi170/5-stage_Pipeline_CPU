/***************************************************
Student Name: 李懿麒 陳品戎
Student ID: 0816032 0816102
***************************************************/

module Hazard_detection(
	input [4:0] IFID_regRs,
	input [4:0] IFID_regRt,
	input [4:0] IDEXE_regRd,
	input IDEXE_memRead,
	output PC_write,
	output IFID_write,
	output control_output_select
);


endmodule

